module notify

pub enum Level {
	low
	normal
	critical
}
